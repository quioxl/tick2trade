`include "uvm_macros.svh"
package system_env_pkg;
  import uvm_pkg::*;
  import avalon_pkg::*;
  import feed_agent_pkg::*;
  import host_agent_pkg::*;
  import order_pkg::*;
  import symbol_map_pkg::*;
  import feed_env_pkg::*;
  import strategy_env_pkg::*;

  //Classes
  `include "system_env_config.svh"
  `include "system_env.svh"
  
endpackage : system_env_pkg
  