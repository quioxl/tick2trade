`include "uvm_macros.svh"
package feed_env_pkg;
  import uvm_pkg::*;
  import avalon_pkg::*;

  `include "feed_message_item.svh"
  `include "feed_message_to_avalon_seq.svh"
  `include "feed_env_config.svh"
  `include "feed_layering.svh"
  `include "feed_env.svh"
  `include "feed_simple_seq.svh"
endpackage