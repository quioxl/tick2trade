`include "uvm_macros.svh"
package system_test_pkg;
  import uvm_pkg::*;
  import avalon_pkg::*;
  import feed_agent_pkg::*;
  import host_agent_pkg::*;
  import order_pkg::*;
  import system_env_pkg::*;
  import strategy_seq_pkg::*;
  import system_seq_pkg::*;

  `include "system_test_base.svh"
  `include "sanity_test.svh"
  //`include "basic_test.svh"
  `include "all_messages_test.svh"
  
endpackage : system_test_pkg
