// ---------------------------------------------------------------------------
//
//  Copyright 2014 IMC. All Rights Reserved.
//
//  Description: Common elements to the Strategy blocks
//
// ---------------------------------------------------------------------------
package strat_pkg;


endpackage