`include "uvm_macros.svh"
package feed_agent_pkg;
  import uvm_pkg::*;
  import avalon_pkg::*;
  `include "feed_message_item.svh"
  `include "feed_message_to_avalon_seq.svh"
  `include "feed_monitor.svh"
  `include "feed_layering.svh"
  `include "feed_simple_seq.svh"
  `include "feed_random_seq.svh"
endpackage