interface order_interface;
  logic clk;
  logic reset_n;
  logic [127:0] data;
  logic ready;
  logic valid;
endinterface