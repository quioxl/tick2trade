// ---------------------------------------------------------------------------
//
//  Copyright 2014 IMC. All Rights Reserved.
//
//  Description: Common elements to the Tick2Trade blocks
//
// ---------------------------------------------------------------------------
package t2t_pkg;

  // Message Type encoding
  parameter  MSG_NEW           = 24'h4E_45_57; // ASCII "NEW"

endpackage
