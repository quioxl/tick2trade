`include "uvm_macros.svh"
package feed_env_pkg;
  import uvm_pkg::*;
  import avalon_pkg::*;

  `include "feed_env_config.svh"
  `include "feed_env.svh"
endpackage