`include "uvm_macros.svh"

package order_out_pkg;
  import uvm_pkg::*;

  `include "order_item.svh";
  `include "order_config.svh";
  `include "order_driver.svh";
  `include "order_monitor.svh"
  `include "order_agent.svh";
endpackage