mhorn@cob-mhorn-centos.4387:1485203932